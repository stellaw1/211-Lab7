module ALU_tb();
    reg [15:0] sim_Ain, sim_Bin;
    reg [1:0] sim_ALUop;
    reg err;
    wire [15:0] sim_out;
    wire sim_Z;


endmodule