module shifter_tb();
    reg [15:0] sim_in;
    reg [1:0] sim_shift;
    reg err;
    wire [15:0] sim_sout;


endmodule