//include finite state machine controller (Controller), an instruction register, an instruction decoder and a datapath
module lab6_top();


endmodule