module regfile_tb();
    reg [15:0] sim_data_in;
    reg [2:0] sim_writenum, sim_readnum;
    reg sim_write, sim_clk;
    reg err;
    wire [15:0] sim_data_out;

    

endmodule