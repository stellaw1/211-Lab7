module datapath(mdata, sximm8, sximm5, vsel, writenum, write, readnum, clk, loada, loadb, loadc, loads, shift, asel, bsel, ALUop, V, N, Z, datapath_out);
    input [15:0] mdata; //16-bit output of a memory block (Lab7)
    input [15:0] sximm8; //sign extended 8-bit immediate driven from instruction decoder. sximm8 is a 16-bit sign extended version of the 8-bit value in the lower 8-bits of the instruction register
    input [15:0] sximm5;
    input write, clk, loada, loadb, loadc, loads, asel, bsel;
    input [3:0] vsel;
    input [2:0] writenum, readnum;
    input [1:0] shift, ALUop;
    output V, N, Z;
    output [15:0] datapath_out;

    //declare signals
    wire[15:0] data_in, data_out, fromAtoMux6, fromBtoShifter, sout, Ain, Bin, out;
    wire[7:0] PC;
    wire [2:0] status;

    //assign zero to mdata and PC
    assign mdata = 16'b0;
    assign PC = 8'b0;

    //instantiate block 9: first 4 bit one-hot MUX. 
    //  vsel = 1000: mdata
    //  vsel = 0100: sximm8
    //  vsel = 0010: {8'b0, PC}
    //  vsel = 0001: datapath_out
    Mux4 #(16) mux1(mdata, sximm8, {8'b0, PC}, datapath_out, vsel, data_in);

    //instantiate block 1: register file
    regfile REGFILE(data_in, writenum, write, readnum, clk, data_out);

    //instantiat blocks 3 and 4: pipeline register A and B
    vDFFE #(16) pipeA(clk, loada, data_out, fromAtoMux6); 
    vDFFE #(16) pipeB(clk, loadb, data_out, fromBtoShifter); 

    //instantiate block 8: shifter unit
    shifter shifter8(fromBtoShifter, shift, sout);  

    //instantiate block 6 and 7: Mux6 and Mux7
    assign Ain = asel ? 16'b0 : fromAtoMux6;
    assign Bin = bsel ? sximm5 : sout;

    //instantiate block 2: ALU unit
    ALU alu2(Ain, Bin, ALUop, out, status); //status[0]=Z, status[1]=N, status[2]=V

    //instantiate block 5: pipeline register C
    vDFFE #(16) pipeC(clk, loadc, out, datapath_out);

    //instantiate block 10: 3-bit status register
    vDFFE #(3) status10(clk, loads, status, {V, N, Z});
endmodule